library IEEE;
Use IEEE.STD_LOGIC_1164.ALL;
USe IEEE.NUMERIC_STD.ALL;

entity rom is
    Generic(
        ADDR_WIDTH : integer:= 7;
        DATA_WIDTH : integer:= 8
    );
    Port ( clk : in STD_LOGIC;
    addr_r: in STD_LOGIC_VECTOR (ADDR_WIDTH-1 downto 0);
     data : out STD_LOGIC_VECTOR (DATA_WIDTH-1 downto 0));
end rom;

Architecture Behavioral of rom is
constant ROM_DEPTH: integer := 2**ADDR_WIDTH-1;   -- but we havent used all of them, only a to as has been used.
type rom_type is array (0 to 98) of std_logic_vector (DATA_WIDTH-1 downto 0);
constant D1_ROM: rom_type :=
(
"00000000",
"00000001",
"00000010",
"00000011",
"00000100",
"00000101",
"00000110",
"00000111",
"00001000",
"00001001",
"00010000",
"00010001",
"00010010",
"00010011",
"00010100",
"00010101",
"00010110",
"00010111",
"00011000",
"00011001",
"00100000",
"00100001",
"00100010",
"00100011",
"00100100",
"00100101",
"00100110",
"00100111",
"00101000",
"00101001",
"00110000",
"00110001",
"00110010",
"00110011",
"00110100",
"00110101",
"00110110",
"00110111",
"00111000",
"00111001",
"01000000",
"01000001",
"01000010",
"01000011",
"01000100",
"01000101",
"01000110",
"01000111",
"01001000",
"01001001",
"01010000",
"01010001",
"01010010",
"01010011",
"01010100",
"01010101",
"01010110",
"01010111",
"01011000",
"01011001",
"01100000",
"01100001",
"01100010",
"01100011",
"01100100",
"01100101",
"01100110",
"01100111",
"01101000",
"01101001",
"01110000",
"01110001",
"01110010",
"01110011",
"01110100",
"01110101",
"01110110",
"01110111",
"01111000",
"01111001",
"10000000",
"10000001",
"10000010",
"10000011",
"10000100",
"10000101",
"10000110",
"10000111",
"10001000",
"10001001",
"10010001",
"10010010",
"10010011",
"10010100",
"10010101",
"10010110",
"10010111",
"10011000",
"10011001"
);

signal rom: rom_type;
begin
    process (clk)
    begin
        if (clk'event and clk = '1') then
            data <= D1_ROM(to_integer(unsigned (addr_r)));
        end if;
    end process;
end Behavioral;